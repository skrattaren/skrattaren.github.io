.. title: Nyårspresenter
.. slug: presenter
.. date: 2007-01-14 15:01:51
.. tags: 

Mitt vild svin i sitt hus. Tack till
`Marria <http://my.opera.com/gagnjungfrun/>`__ och
`Dinara <http://my.opera.com/trolljomfru/>`__!


(-%E

|image0|

.. |image0| image:: http://files.myopera.com/Sterkrig/blog/svin_i_sitt_hus.jpg
