.. title: Ásmegin: fotto
.. slug: asmegin-fotto
.. date: 2007-02-05 20:02:37
.. tags: sve,musik,рус,eng

Ásmegins fotografialbum om inspelning av det nya CD:

`Ásmegin <http://www.asmegin.com/Galleri/index.php?gallery=Recordings%20of%20the%20new%20album>`__
