.. title: "sterkrig"
.. slug: sterkrig-is-min-nama
.. date: 2007-04-01 17:04:38
.. tags: sve,рус,eng

Jag har ett riktigt svenskt namn (-:E Google har funnit endast
`pdf-filen <http://www.vasttrafik.se/directory/publications/51188/Pling%20060908.pdf>`__
inte om mig själv 4-:E
