.. title: Font
.. slug: font
.. date: 2007-03-19 22:03:56
.. tags: 

Vem vet vad teckesnitt är det?

|image0|

.. |image0| image:: http://files.myopera.com/Sterkrig/blog/teckensnitt.png
