.. title: Nils Olav III den norsk ridder
.. slug: den-norsk-ridder
.. date: 2008-08-20 12:08:47
.. tags: sve,рус,linux,eng

|image0|

Kungspingvin Nils Olav III har blivit en norsk riddare och överste av
Hans Majestet Kongens Garde

`Läs på norska...
<http://www.vg.no/nyheter/utrolige-historier/artikkel.php?artid=524663>`__

`Mer... <http://www.nrk.no/nyheter/utenriks/1.6178426>`__

Schelmish - Igni Gena (2004)

.. |image0| image:: http://www.nrk.no/contentfile/file/1.6178592!f169CropList/img650x367.jpg
