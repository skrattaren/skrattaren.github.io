.. title: IMified
.. slug: imified
.. date: 2007-10-28 00:10:45
.. tags: sve,рус,eng,jabber

Jag kunde skriva om `IMified <http://imified.com/>`__, därför att det
verkar slutligen... Men du skall hellre läsa om det på dess huvudsiden i
engelska, du kan, tror jag (-;E

Och dessa engelska skulle våra förståeligare för alla än min
svenska…
