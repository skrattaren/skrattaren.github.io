.. title: Íslenska
.. slug: islenska
.. date: 2006-12-17 17:12:18
.. tags: lang

Есть в древнеисландском хорошее слово — **hraustr**. И значит оно
*"доблестный, сильный"*. Красивое слово, звучное. Считается, что
восходит к общеиндоевропейскому корню. И в русском языке этот корень
представлен словом **"крот"**.

У древних германцев и древних славян представления о доблести и силе
определённо несколько расходились (-%Е

-------------

There's a good word in Old Icelandic, **hraustr** (meaning *brave,
strong*). Sounds conformably. It's believed to be derived from
Indoeuropean root, and this root is presented in Russian as **"крот"**
(*[krot]*, a mole)

Ancient Teutons and Slavs seem to me to have a little bit different
conception of strength and valour (-%E

-------------

Det finns ett gott ord i fornisländska — **hraustr**. Det betyder
*kraftig, modig, djärv*. Och ljuder det lika så. Detta ord är trott att
härstamma från Indoeuropiska språket, och dessa ordrot finns i Ryska, i
ett ord **"крот"** (*[krot]*, mullvad)

Fornslaver och -germaner föreväller hava en lite skild föreställning
om kraft o s v (-%E
