.. title: Edicode
.. slug: edicode
.. date: 2006-12-07 16:12:08
.. tags: 

Показал мне как-то `**LoiR** <http://my.opera.com/LoiR/about/>`__ `вот
такую
штуку <http://www.guntherkrauss.de/computer/xml/daten/edicode.html>`__ —
панельку с всякими раскрасивыми unicode-символами. Добавляем себе в
боковую панель и радуемся удобной вставке символов, коды которых не
упомнить (-:Е

About two weeks ago `**LoiR** <http://my.opera.com/LoiR/about/>`__, a
friend of mine, pointed
`Edicode <http://www.guntherkrauss.de/computer/xml/daten/edicode.html>`__
sidebar out for me. If you have to deal with non-ASCII symbols, absent
in your keyboard layout, then that's tool you need (-:E

`**LoiR** <http://my.opera.com/LoiR/about/>`__ den vännen min visade mig
`Edicode
sidpanelen <http://www.guntherkrauss.de/computer/xml/daten/edicode.html>`__.
Nu kan jag klistra var unicode-tecken som jag behöver in (-:E

Hagalaz' Runedance - The Winds That Sang Of Midgard's Fate [1998]
