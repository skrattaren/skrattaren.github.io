.. title: Den krigaren av Öppna Källkod
.. slug: OK-krigaren
.. date: 2007-10-19 15:10:00
.. tags: sve,рус,linux,eng

Jag är den store krigaren av Öppna Källkod! Kubuntu_ och Xubuntu_ 7.10 vår
utgivat igår och på densamma kväll har jag alla åtta CD-avbilder av Kubuntu och
Xubuntu nedladdat och framlagt dem i lokalnätverk, för alla att försöka eller
installera. Och idag jag laddade två avbilder upp för Ubuntu-användare ute i
Fjärran Öst (-:E

.. _Kubuntu: http://kubuntu.org/announcements/7.10-release.php
.. _Xubuntu: http://xubuntu.org/news/gutsy/release

Веснянка - Ой, заграли музиченьки [2003]
