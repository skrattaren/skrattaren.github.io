.. title: digiKam: Menyrad
.. slug: digikam-menyrad
.. date: 2008-01-04 22:01:06
.. tags: sve,рус,linux,eng

Vill du möjliggöra menyrad i `digiKam <http://www.digikam.org/>`__? Se
här!


 ***sterkrig@trollsdatorn ~ $** nano ~/.kde/share/config/digikamrc*

::

    [MainWindow]

    MenuBar=Enabled

