.. title: Bandbrytande nyheter!
.. slug: nyheter
.. date: 2007-05-16 01:05:58
.. tags: sve,рус,eng,хе-хе

    The Orthoptera are the only insects considered kosher in Judaism


(***Wikipedia***)
